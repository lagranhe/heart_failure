�csklearn.ensemble._forest
RandomForestClassifier
q )�q}q(X   base_estimatorqcsklearn.tree._classes
DecisionTreeClassifier
q)�q}q(X	   criterionqX   giniqX   splitterq	X   bestq
X	   max_depthqNX   min_samples_splitqKX   min_samples_leafqKX   min_weight_fraction_leafqG        X   max_featuresqNX   max_leaf_nodesqNX   random_stateqNX   min_impurity_decreaseqG        X   class_weightqNX	   ccp_alphaqG        X   _sklearn_versionqX   1.0.1qubX   n_estimatorsqKX   estimator_paramsq(hhhhhhhhhhtqX	   bootstrapq�X	   oob_scoreq�X   n_jobsqNhK X   verboseqK X
   warm_startq�hNX   max_samplesqNhhhNhKhKhG        hX   autoq hNhG        hG        X   feature_names_in_q!cnumpy.core.multiarray
_reconstruct
q"cnumpy
ndarray
q#K �q$Cbq%�q&Rq'(KK�q(cnumpy
dtype
q)X   O8q*���q+Rq,(KX   |q-NNNJ����J����K?tq.b�]q/(X   ageq0X   anaemiaq1X   creatinine_phosphokinaseq2X   diabetesq3X   ejection_fractionq4X   high_blood_pressureq5X	   plateletsq6X   serum_creatinineq7X   serum_sodiumq8X   sexq9X   smokingq:etq;bX   n_features_in_q<KX
   n_outputs_q=KX   classes_q>h"h#K �q?h%�q@RqA(KK�qBh)X   i8qC���qDRqE(KX   <qFNNNJ����J����K tqGb�C               qHtqIbX
   n_classes_qJKX   base_estimator_qKhX   estimators_qL]qM(h)�qN}qO(hhh	h
hNhKhKhG        hh hNhJ�
hG        hNhG        h<Kh=Kh>h"h#K �qPh%�qQRqR(KK�qSh)X   f8qT���qURqV(KhFNNNJ����J����K tqWb�C              �?qXtqYbhJcnumpy.core.multiarray
scalar
qZhEC       q[�q\Rq]X   max_features_q^KX   tree_q_csklearn.tree._tree
Tree
q`Kh"h#K �qah%�qbRqc(KK�qdhE�C       qetqfbK�qgRqh}qi(hKX
   node_countqjKSX   nodesqkh"h#K �qlh%�qmRqn(KKS�qoh)X   V56qp���qqRqr(Kh-N(X
   left_childqsX   right_childqtX   featurequX	   thresholdqvX   impurityqwX   n_node_samplesqxX   weighted_n_node_samplesqytqz}q{(hsh)X   i8q|���q}Rq~(KhFNNNJ����J����K tqbK �q�hth~K�q�huh~K�q�hvhVK�q�hwhVK �q�hxh~K(�q�hyhVK0�q�uK8KKtq�b�B(         H                    �R@rWW)2��?�             j@       /                  �pAL�9�W�?s             f@                          0`@z�G�z�?U            @_@������������������������       �                     @       *                 l/A@�r-��?P            �]@                          �6@b����o�?6            �R@������������������������       �                     @       !                   �a@b�h�d.�?3            �Q@	                        ����?�?�P�a�?+             N@
                          �F@      �?              @������������������������       �                     �?������������������������       �                     �?                           ��@ܷ��?��?)             M@              	             �?x�}b~|�?(            �L@                            Q@�J�4�?             9@                          �`@���}<S�?             7@������������������������       �                     �?                        pff�?���7�?             6@������������������������       �        
             4@                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @              
             �?      �?             @@������������������������       �                     2@                           �?@4և���?             ,@������������������������       �        	             $@                        ����?      �?             @������������������������       �                      @                          0a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?"       )                   �a@      �?             $@#       (                  x�A����X�?             @$       %                 �p=�?r�q��?             @������������������������       �                     @&       '                    �Q@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @+       ,                   �a@ qP��B�?            �E@������������������������       �                    �C@-       .                   @@@      �?             @������������������������       �                     �?������������������������       �                     @0       5                 `ff�?Np�����?            �I@1       4                 ����?�IєX�?             1@2       3       	             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        
             .@6       C       
             �?�������?             A@7       8                   �;@V�a�� �?             =@������������������������       �                     &@9       >                 ����?�q�q�?	             2@:       ;                    a@      �?              @������������������������       �                     @<       =                   `a@      �?              @������������������������       �                     �?������������������������       �                     �??       B                  XUP@      �?             $@@       A                   �C@����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @D       E                    �I@���Q��?             @������������������������       �                     �?F       G                    �?      �?             @������������������������       �                     @������������������������       �                     �?I       R                   ̊@"pc�
�?            �@@J       O                  @�A     ��?             @@K       N                  @A�>����?             ;@L       M                   a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     8@P       Q                    �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?q�tq�bX   valuesq�h"h#K �q�h%�q�Rq�(KKSKK�q�hV�B0       ``@     �S@     @_@     �I@      Y@      9@              @      Y@      2@      M@      1@              @      M@      (@     �J@      @      �?      �?      �?                      �?      J@      @      J@      @      5@      @      5@       @              �?      5@      �?      4@              �?      �?              �?      �?                       @      ?@      �?      2@              *@      �?      $@              @      �?       @              �?      �?      �?                      �?              �?      @      @       @      @      �?      @              @      �?      �?              �?      �?              �?              @              E@      �?     �C@              @      �?              �?      @              9@      :@      0@      �?      �?      �?      �?                      �?      .@              "@      9@      @      7@              &@      @      (@      �?      @              @      �?      �?      �?                      �?      @      @       @      @              @       @              @              @       @              �?      @      �?      @                      �?      @      ;@      @      ;@       @      9@       @      �?       @                      �?              8@      @       @               @      @              �?        q�tq�bubhhubh)�q�}q�(hhh	h
hNhKhKhG        hh hNhJ/��hG        hNhG        h<Kh=Kh>h"h#K �q�h%�q�Rq�(KK�q�hV�C              �?q�tq�bhJhZhEC       q��q�Rq�h^Kh_h`Kh"h#K �q�h%�q�Rq�(KK�q�hE�C       q�tq�bK�q�Rq�}q�(hKhjKShkh"h#K �q�h%�q�Rq�(KKS�q�hr�B(         D                 p=
�?�=����?�             j@       A                    �T@�W��/�?p            @e@                          �;@ {��e�?k            �c@                          �1@���Q��?             >@������������������������       �                     @       	                    @M@�q�����?             9@                          l�@r�q��?             @������������������������       �                     @������������������������       �                     �?
                          �a@p�ݯ��?             3@                         ��A�t����?             1@                        ����?�C��2(�?             &@������������������������       �                     "@                         ��A      �?              @������������������������       �                     �?������������������������       �                     �?                          Pa@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @       "                   a@X�EQ]N�?V             `@                          @@@d}h���?             E@                         `�A�eP*L��?             &@                           �?      �?              @������������������������       �                     @������������������������       �                      @������������������������       �                     @       !                   ��@��� ��?             ?@                         ��A 	��p�?             =@������������������������       �                     7@                          0�A�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @#       >                     S@ 	��p�?8            �U@$       '                 ����?�IєX�?6            @U@%       &                    �?      �?              @������������������������       �                     �?������������������������       �                     �?(       /                   @@@��`qM|�?4            �T@)       .                    �?�����H�?             "@*       +                   `a@؇���X�?             @������������������������       �                     @,       -                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @0       9                   ;AxL��N�?/            �R@1       2       	             �?"pc�
�?	             &@������������������������       �                     �?3       4                    �?ףp=
�?             $@������������������������       �                     @5       8                   �@      �?             @6       7                  �hA      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @:       =                   �e@ ������?&            �O@;       <                   �c@`2U0*��?             9@������������������������       �                     8@������������������������       �                     �?������������������������       �                     C@?       @                  ��A      �?              @������������������������       �                     �?������������������������       �                     �?B       C                    �?�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?E       J                   �`@��Sݭg�?            �C@F       G                 ���@���N8�?             5@������������������������       �                     3@H       I                    D@      �?              @������������������������       �                     �?������������������������       �                     �?K       P                    �?      �?	             2@L       O                  ��	A      �?              @M       N                   �u@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @Q       R                   ȡ@�z�G��?             $@������������������������       �                     @������������������������       �                     @q�tq�bh�h"h#K �q�h%�q�Rq�(KKSKK�q�hV�B0        a@      R@     �_@     �E@     �_@     �@@      (@      2@              @      (@      *@      @      �?      @                      �?      @      (@      @      (@      �?      $@              "@      �?      �?      �?                      �?      @       @      @                       @       @             �\@      .@     �@@      "@      @      @      @       @      @                       @              @      ;@      @      ;@       @      7@              @       @               @      @                       @     @T@      @      T@      @      �?      �?              �?      �?             �S@      @       @      �?      @      �?      @              @      �?              �?      @               @             �Q@      @      "@       @              �?      "@      �?      @              @      �?      �?      �?      �?                      �?       @              O@      �?      8@      �?      8@                      �?      C@              �?      �?              �?      �?              �?      $@              $@      �?              $@      =@      �?      4@              3@      �?      �?              �?      �?              "@      "@      @       @       @       @               @       @              @              @      @              @      @        q�tq�bubhhubh)�q�}q�(hhh	h
hNhKhKhG        hh hNhJu�7hG        hNhG        h<Kh=Kh>h"h#K �q�h%�q�Rq�(KK�q�hV�C              �?q�tq�bhJhZhEC       q��q�Rq�h^Kh_h`Kh"h#K �q�h%�q�Rq�(KK�q�hE�C       q�tq�bK�q�Rq�}q�(hK	hjKIhkh"h#K �q�h%�q�Rq�(KKI�q�hr�B�         8                 p=
�?�oUN�1�?�             j@                           �?$Z9��?r            �d@              
             �?������?@            @X@                        ����?��ɉ�?+            @P@������������������������       �                    �B@       	                   @@@@4և���?             <@                          ��@z�G�z�?             @������������������������       �                     @������������������������       �                     �?
                         ��@�nkK�?             7@������������������������       �                     6@������������������������       �                     �?                           �T@     ��?             @@                           �N@d}h���?             <@                           �?��S�ۿ?             .@������������������������       �                     $@                          @a@z�G�z�?             @                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @                          �j@�n_Y�K�?             *@������������������������       �                     @                           �?X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                     @       3                   l�@">�֕�?2            �Q@       ,                    �P@b�2�tk�?(             K@       '                 ����?�������?             A@       &                   H�@�>4և��?             <@        !                    �?ȵHPS!�?             :@������������������������       �                     ,@"       %                   �C@      �?
             (@#       $                    �M@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                      @(       )                    �?�q�q�?             @������������������������       �                     @*       +                   �`@�q�q�?             @������������������������       �                     �?������������������������       �                      @-       .                   �`@���Q��?             4@������������������������       �                     @/       2                  `ZA؇���X�?             ,@0       1                   �6@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     $@4       7                    �?      �?
             0@5       6                   �a@�8��8��?             (@������������������������       �                     &@������������������������       �                     �?������������������������       �                     @9       H                   �G@����X�?             E@:       =                   0`@r�q��?             B@;       <                    \@      �?             @������������������������       �                     @������������������������       �                     �?>       G                   ȡ@     ��?             @@?       D                    a@`Jj��?             ?@@       A                 ���@h�����?             <@������������������������       �                     9@B       C                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @E       F                    @P@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @q�tq�bh�h"h#K �q�h%�q�Rq�(KKIKK�q�hV�B�        b@      P@     �`@      A@     @U@      (@     �O@       @     �B@              :@       @      @      �?      @                      �?      6@      �?      6@                      �?      6@      $@      6@      @      ,@      �?      $@              @      �?       @      �?       @                      �?       @               @      @      @              @      @      @                      @              @      H@      6@     �@@      5@      9@      "@      7@      @      7@      @      ,@              "@      @      @      @              @      @              @                       @       @      @              @       @      �?              �?       @               @      (@      @               @      (@       @       @               @       @                      $@      .@      �?      &@      �?      &@                      �?      @              (@      >@      @      >@      @      �?      @                      �?      @      =@       @      =@      �?      ;@              9@      �?       @      �?                       @      �?       @               @      �?              �?              @        q�tq�bubhhubh)�q�}q�(hhh	h
hNhKhKhG        hh hNhJ��!XhG        hNhG        h<Kh=Kh>h"h#K �q�h%�q�Rq�(KK�q�hV�C              �?q�tq�bhJhZhEC       qنq�Rq�h^Kh_h`Kh"h#K �q�h%�q�Rq�(KK�q�hE�C       q�tq�bK�q�Rq�}q�(hK	hjKOhkh"h#K �q�h%�q�Rq�(KKO�q�hr�BH                            �`@��+s�?�             j@                          0�@���Q��?'             N@                          �`@����X�?            �H@                          �P@H%u��?             9@                          �B@      �?              @������������������������       �                     �?������������������������       �                     �?                          A���}<S�?             7@	       
                    @F@���7�?             6@������������������������       �                     �?������������������������       �                     5@������������������������       �                     �?                          �C@r�q��?             8@                           �R@���Q��?             4@                        p=
�?���!pc�?             &@������������������������       �                      @������������������������       �                     @������������������������       �                     "@                           �?      �?             @������������������������       �                     @������������������������       �                     �?                          ��@�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?       &                  ��	A�Ҳ���?^            �b@                        pff�?      �?             <@                           �?d}h���?             ,@������������������������       �                      @                          H�@      �?             @������������������������       �                     @������������������������       �                     @        !                   �@d}h���?	             ,@������������������������       �                     "@"       #                  �CA���Q��?             @������������������������       �                      @$       %                    �Q@�q�q�?             @������������������������       �                     �?������������������������       �                      @'       N                   ʶ@�)l�o��?J            @^@(       ;                   @@@p�5�9��?I            �]@)       ,                    �I@��S���?             >@*       +                   Ж@      �?              @������������������������       �                     @������������������������       �                     �?-       2                    �?�X����?             6@.       1                    �P@z�G�z�?             $@/       0                   �w@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @3       6                 ����?�q�q�?             (@4       5                   @a@r�q��?             @������������������������       �                     �?������������������������       �                     @7       :                   �a@�q�q�?             @8       9       	             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @<       E                    �?������?4            @V@=       D                   `e@ 7���B�?             K@>       C                   �b@�����?             5@?       @                   �K@P���Q�?             4@������������������������       �                     1@A       B                   �^@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                    �@@F       G                   A؇���X�?            �A@������������������������       �                     :@H       M                    �?X�<ݚ�?             "@I       L       
             �?�q�q�?             @J       K                  �W A�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @q�tq�bh�h"h#K �q�h%�q�Rq�(KKOKK�q�hV�B�       �`@     �R@      8@      B@      ,@     �A@      @      6@      �?      �?      �?                      �?       @      5@      �?      5@      �?                      5@      �?              &@      *@       @      (@       @      @       @                      @              "@      @      �?      @                      �?      $@      �?      $@                      �?     �[@     �C@      ,@      ,@      &@      @       @              @      @      @                      @      @      &@              "@      @       @       @              �?       @      �?                       @      X@      9@      X@      7@      ,@      0@      @      �?      @                      �?      @      .@       @       @       @      @              @       @                      @      @      @      �?      @      �?                      @      @       @      �?       @               @      �?              @             �T@      @      J@       @      3@       @      3@      �?      1@               @      �?       @                      �?              �?     �@@              >@      @      :@              @      @      @       @      �?       @               @      �?              @                      @               @q�tq�bubhhubh)�q�}q�(hhh	h
hNhKhKhG        hh hNhJC�NhG        hNhG        h<Kh=Kh>h"h#K �q�h%�q�Rq�(KK�q�hV�C              �?q�tq�bhJhZhEC       q��q�Rq�h^Kh_h`Kh"h#K �q�h%�q�Rq�(KK�q�hE�C       r   tr  bK�r  Rr  }r  (hKhjKQhkh"h#K �r  h%�r  Rr  (KKQ�r  hr�B�         @                    �R@⚥?��?�             j@                          0`@�h{���?o            `f@                            F@�t����?             1@������������������������       �                     @                          ��@؇���X�?             ,@������������������������       �                     (@������������������������       �                      @                          �;@�{��?��?g            @d@	                           @L@��}*_��?             ;@
                         �?A8�Z$���?             *@                         �2A���Q��?             @������������������������       �                      @              
             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @                          pi@և���X�?	             ,@                          �`@؇���X�?             @������������������������       �                     @                            O@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @       9                   ��@�T�H���?W            �`@       2                     @����y7�?R            @_@       /       	             �?io8�?K             ]@       .       
             �?R���Q�?             D@                           �H@�ݜ�?            �C@������������������������       �        	             *@       -                   ؂@���B���?             :@                         pff�?�E��ӭ�?             2@������������������������       �                     �?!       (                     Q@������?             1@"       '                   �|@؇���X�?
             ,@#       $                   pa@$�q-�?	             *@������������������������       �                     "@%       &                  0�A      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?)       *                   �`@�q�q�?             @������������������������       �                     �?+       ,                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?0       1                 ����?�"w����?-             S@������������������������       �                     �?������������������������       �        ,            �R@3       6       
             �?X�<ݚ�?             "@4       5                   �F@      �?             @������������������������       �                     @������������������������       �                     �?7       8                 ���@���Q��?             @������������������������       �                      @������������������������       �                     @:       ?                  ��A���Q��?             $@;       <                    @H@և���X�?             @������������������������       �                     @=       >                 LXA      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @A       P                   (�@������?             >@B       G                   �D@�+$�jP�?             ;@C       D                   �`@�IєX�?             1@������������������������       �                     &@E       F                   a@r�q��?             @������������������������       �                     �?������������������������       �                     @H       O       
             �?���Q��?             $@I       N                   �K@և���X�?             @J       K                  8�A���Q��?             @������������������������       �                      @L       M                   �r@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     @r	  tr
  bh�h"h#K �r  h%�r  Rr  (KKQKK�r  hV�B       �a@     �P@     �`@     �F@      @      (@      @               @      (@              (@       @              `@     �@@      $@      1@       @      &@       @      @               @       @      �?       @                      �?               @       @      @      �?      @              @      �?       @               @      �?              @             �]@      0@     @\@      (@     @[@      @      A@      @      A@      @      *@              5@      @      *@      @              �?      *@      @      (@       @      (@      �?      "@              @      �?      @                      �?              �?      �?       @              �?      �?      �?              �?      �?               @                      �?     �R@      �?              �?     �R@              @      @      �?      @              @      �?              @       @               @      @              @      @      @      @              @      @      �?              �?      @              @               @      6@      @      6@      �?      0@              &@      �?      @      �?                      @      @      @      @      @       @      @               @       @      �?              �?       @               @                      @      @        r  tr  bubhhubh)�r  }r  (hhh	h
hNhKhKhG        hh hNhJ�R�[hG        hNhG        h<Kh=Kh>h"h#K �r  h%�r  Rr  (KK�r  hV�C              �?r  tr  bhJhZhEC       r  �r  Rr  h^Kh_h`Kh"h#K �r  h%�r  Rr  (KK�r  hE�C       r   tr!  bK�r"  Rr#  }r$  (hK
hjKMhkh"h#K �r%  h%�r&  Rr'  (KKM�r(  hr�B�         >                 p=
�?Z��s�N�?�             j@       !                    �?,zmYA��?l            �e@                           *�@\������?>            @Z@                          �`@�+e�X�?:             Y@                           �?      �?	             0@������������������������       �                     @                         8�Ar�q��?             (@������������������������       �                     @	       
                     S@�q�q�?             @������������������������       �                      @������������������������       �                     @                           �?r�q��?1             U@������������������������       �                     F@                          @@@��Q��?             D@                          �a@������?	             .@                          �;@d}h���?             ,@������������������������       �                      @                           b@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     �?                           �Q@H%u��?             9@                          �K@���7�?             6@������������������������       �        
             1@                           �?z�G�z�?             @������������������������       �                      @                          �x@�q�q�?             @������������������������       �                      @������������������������       �                     �?              
             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @"       =                   �@H�V�e��?.             Q@#       ,                     K@p�v>��?!            �G@$       )                  ��A      �?             2@%       (       	             �?�q�q�?             (@&       '                    �?�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @*       +                    �H@r�q��?             @������������������������       �                     �?������������������������       �                     @-       8                   @@@д>��C�?             =@.       /                 ����?և���X�?             @������������������������       �                     �?0       1                    �?�q�q�?             @������������������������       �                      @2       3                 ����?      �?             @������������������������       �                     �?4       5                   �`@�q�q�?             @������������������������       �                     �?6       7                   a@      �?              @������������������������       �                     �?������������������������       �                     �?9       <                   �`@���7�?             6@:       ;       	             �?؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     .@������������������������       �                     5@?       @                  ���@�E��ӭ�?             B@������������������������       �                     @A       F                   �`@�'�`d�?            �@@B       C                   0�@���7�?             6@������������������������       �                     3@D       E                 Уp�?�q�q�?             @������������������������       �                      @������������������������       �                     �?G       H                 ��� @�eP*L��?             &@������������������������       �                     @I       L       	             �?      �?              @J       K                  ��A      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @r)  tr*  bh�h"h#K �r+  h%�r,  Rr-  (KKMKK�r.  hV�B�       �a@     @Q@     @`@     �E@      S@      =@      S@      8@      @      $@      @               @      $@              @       @      @       @                      @     �Q@      ,@      F@              :@      ,@      @      &@      @      &@               @      @      @              @      @              �?              6@      @      5@      �?      1@              @      �?       @               @      �?       @                      �?      �?       @               @      �?                      @      K@      ,@     �@@      ,@      "@      "@       @      @       @      @       @                      @      @              �?      @      �?                      @      8@      @      @      @      �?               @      @               @       @       @              �?       @      �?      �?              �?      �?              �?      �?              5@      �?      @      �?              �?      @              .@              5@              $@      :@      @              @      :@      �?      5@              3@      �?       @               @      �?              @      @              @      @       @       @       @       @                       @      @        r/  tr0  bubhhubh)�r1  }r2  (hhh	h
hNhKhKhG        hh hNhJ�v}hG        hNhG        h<Kh=Kh>h"h#K �r3  h%�r4  Rr5  (KK�r6  hV�C              �?r7  tr8  bhJhZhEC       r9  �r:  Rr;  h^Kh_h`Kh"h#K �r<  h%�r=  Rr>  (KK�r?  hE�C       r@  trA  bK�rB  RrC  }rD  (hK
hjK_hkh"h#K �rE  h%�rF  RrG  (KK_�rH  hr�B�         "                   �`@⚥?��?�             j@                           �R@<��¤�?'             Q@                          �6@v ��?            �E@                           @J@      �?              @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @	                        ����?<=�,S��?            �A@
                         ��Ar�q��?             2@������������������������       �                     �?              	             �?�t����?             1@                          �a@      �?              @������������������������       �                     �?                          �v@؇���X�?             @                          �l@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@              	             �?j���� �?             1@������������������������       �                     @                          �`@�z�G��?             $@                           �?      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                      @                        ����?�J�4�?             9@������������������������       �                      @                           �T@���}<S�?             7@������������������������       �                     *@        !                   P�@z�G�z�?             $@������������������������       �                      @������������������������       �                      @#       X                     S@:��o#@�?^            �a@$       M                    �P@�����?X            �`@%       :                  ��A�?�'�@�?I            �\@&       -                    �?,�+�C�?"            �K@'       (                   Pa@z�G�z�?             $@������������������������       �                     @)       ,                    �?���Q��?             @*       +                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @.       /                 ����?`Ӹ����?            �F@������������������������       �                     6@0       3       	             �?���}<S�?             7@1       2                   �}@�q�q�?             @������������������������       �                      @������������������������       �                     �?4       9                   �;@P���Q�?             4@5       8                  ��	A؇���X�?             @6       7                   0a@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     *@;       >                    �?F�4�Dj�?'            �M@<       =                  ��@�7��?            �C@������������������������       �                    �B@������������������������       �                      @?       @                   a@�G�z��?             4@������������������������       �                     @A       H                   @s@ҳ�wY;�?             1@B       G                   pg@X�<ݚ�?             "@C       F                    �?z�G�z�?             @D       E                 033�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @I       L                    �?      �?              @J       K                   ��@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @N       S                    �?�z�G��?             4@O       P                 p=
�?8�Z$���?	             *@������������������������       �                     "@Q       R                   0a@      �?             @������������������������       �                      @������������������������       �                      @T       U                    >@և���X�?             @������������������������       �                     @V       W                    I@      �?             @������������������������       �                     @������������������������       �                     �?Y       ^                   @J@����X�?             @Z       ]                 ����?r�q��?             @[       \                   @a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?rI  trJ  bh�h"h#K �rK  h%�rL  RrM  (KK_KK�rN  hV�B�       �a@     �P@      ;@     �D@      7@      4@      �?      @      �?      �?              �?      �?                      @      6@      *@      .@      @              �?      .@       @      @       @              �?      @      �?       @      �?       @                      �?      @              "@              @      $@              @      @      @      @      �?              �?      @                       @      @      5@       @               @      5@              *@       @       @               @       @             �\@      :@     @\@      5@     �X@      .@     �I@      @       @       @      @              @       @      �?       @      �?                       @       @             �E@       @      6@              5@       @       @      �?       @                      �?      3@      �?      @      �?       @      �?              �?       @              @              *@              H@      &@     �B@       @     �B@                       @      &@      "@              @      &@      @      @      @      @      �?      �?      �?      �?                      �?      @                      @      @      �?      @      �?      @                      �?      @              ,@      @      &@       @      "@               @       @       @                       @      @      @              @      @      �?      @                      �?       @      @      �?      @      �?      �?      �?                      �?              @      �?        rO  trP  bubhhubh)�rQ  }rR  (hhh	h
hNhKhKhG        hh hNhJg}�XhG        hNhG        h<Kh=Kh>h"h#K �rS  h%�rT  RrU  (KK�rV  hV�C              �?rW  trX  bhJhZhEC       rY  �rZ  Rr[  h^Kh_h`Kh"h#K �r\  h%�r]  Rr^  (KK�r_  hE�C       r`  tra  bK�rb  Rrc  }rd  (hKhjKahkh"h#K �re  h%�rf  Rrg  (KKa�rh  hr�B8         $                   �`@
��P ��?�             j@                          �C@�d�����?/            @R@                           `S@��i#[�?             E@                          �U@<=�,S��?            �A@������������������������       �                     @                        p=
�?�P�*�?             ?@                          RAև���X�?             5@       	                   p`@      �?              @������������������������       �                     @
                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?              	             �?�θ�?             *@                         �?Aև���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @                          �`@ףp=
�?	             $@������������������������       �                      @                            P@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                          �Af���M�?             ?@������������������������       �                     @                        `ff�?����X�?             <@������������������������       �                     @       #                    �?�ՙ/�?             5@                         �Aև���X�?             ,@������������������������       �                      @                            �?�q�q�?             (@������������������������       �                     @!       "                   Xt@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     @%       8                   �;@��¤��?_             a@&       -                   Pa@և���X�?             <@'       (                  ��	A�q�q�?             (@������������������������       �                     @)       *                    �?�����H�?             "@������������������������       �                     @+       ,                   a@�q�q�?             @������������������������       �                     �?������������������������       �                      @.       1                   �a@      �?             0@/       0                 ����?�����H�?             "@������������������������       �                      @������������������������       �                     �?2       5                    �?և���X�?             @3       4       	             �?      �?             @������������������������       �                     @������������������������       �                     �?6       7                   Hr@�q�q�?             @������������������������       �                     �?������������������������       �                      @9       Z                   �L@4?,R��?L             [@:       K                  pA��l��?C            @X@;       J                  ��@xdQ�m��?7            @T@<       =                   @B@P���Q�?6             T@������������������������       �                     @@>       I                    �U@�8��8��?              H@?       F                    �?�nkK�?             G@@       E                   @a@`���i��?             F@A       B                 �uA�8��8��?             (@������������������������       �                     "@C       D                   �C@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @@G       H                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?L       O                 `ff�?      �?             0@M       N                  poA؇���X�?             @������������������������       �                     @������������������������       �                     �?P       U                    �J@X�<ݚ�?             "@Q       T       
             �?      �?             @R       S       	             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @V       W       
             �?z�G�z�?             @������������������������       �                     @X       Y                 pff�?      �?              @������������������������       �                     �?������������������������       �                     �?[       `                    �?���|���?	             &@\       _       	             �?      �?              @]       ^                   ��@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @ri  trj  bh�h"h#K �rk  h%�rl  Rrm  (KKaKK�rn  hV�B       @a@     �Q@     �@@      D@      *@      =@      *@      6@              @      *@      2@      (@      "@       @      @              @       @      �?       @                      �?      $@      @      @      @      @                      @      @              �?      "@               @      �?      �?      �?                      �?              @      4@      &@              @      4@       @      @              *@       @      @       @       @              @       @              @      @      @              @      @              @             @Z@      ?@      (@      0@       @      @              @       @      �?      @               @      �?              �?       @              @      (@      �?       @               @      �?              @      @      �?      @              @      �?               @      �?              �?       @             @W@      .@     �U@      &@      S@      @      S@      @      @@              F@      @      F@       @     �E@      �?      &@      �?      "@               @      �?              �?       @              @@              �?      �?      �?                      �?               @              �?      $@      @      @      �?      @                      �?      @      @      @      �?      �?      �?      �?                      �?       @              �?      @              @      �?      �?      �?                      �?      @      @      @      @      �?      @              @      �?              @              @        ro  trp  bubhhubh)�rq  }rr  (hhh	h
hNhKhKhG        hh hNhJ	�tlhG        hNhG        h<Kh=Kh>h"h#K �rs  h%�rt  Rru  (KK�rv  hV�C              �?rw  trx  bhJhZhEC       ry  �rz  Rr{  h^Kh_h`Kh"h#K �r|  h%�r}  Rr~  (KK�r  hE�C       r�  tr�  bK�r�  Rr�  }r�  (hK	hjKGhkh"h#K �r�  h%�r�  Rr�  (KKG�r�  hr�B�         $                   �q@V2�d��?�             j@                        p=
�?hb�Iy��?@            @[@                           �T@���X�?"             L@                          �;@��x_F-�?             �I@������������������������       �                     @                         �wA�q��/��?             G@                           n@ �#�Ѵ�?            �E@       	                  �A�Ń��̧?             E@������������������������       �                     C@
              
             �?      �?             @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @                          `c@䯦s#�?            �J@                         �m
A�E��ӭ�?             B@������������������������       �                     (@                            R@�q�q�?             8@                           �?���Q��?             .@������������������������       �                     @                           �?�q�q�?             "@������������������������       �                     @������������������������       �                     @                           a@�����H�?             "@������������������������       �                      @������������������������       �                     �?       #                    m@j���� �?	             1@       "                   �f@�θ�?             *@        !                    d@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @%       F                   <�@z�G�z�?B             Y@&       7                  �Ar�q��??             X@'       ,                   �`@�eP*L��?             6@(       )                   �C@      �?              @������������������������       �                     @*       +                    @I@�q�q�?             @������������������������       �                      @������������������������       �                     �?-       0                   �@d}h���?             ,@.       /                    �?      �?              @������������������������       �                     �?������������������������       �                     �?1       2                   �a@r�q��?             (@������������������������       �                     @3       6                    �?���Q��?             @4       5                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @8       A                    �?�L���?-            �R@9       @                   ��@z�G�z�?             9@:       ;                    �Q@      �?             4@������������������������       �                     ,@<       ?                    `S@r�q��?             @=       >                   �B@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @B       C                 p=
�?@�E�x�?            �H@������������������������       �                    �F@D       E                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KKGKK�r�  hV�Bp       �a@      Q@     �N@      H@     �D@      .@     �D@      $@              @     �D@      @     �D@       @     �D@      �?      C@              @      �?      �?      �?      �?                      �?       @                      �?              @              @      4@     �@@      $@      :@              (@      $@      ,@      "@      @      @              @      @      @                      @      �?       @               @      �?              $@      @      $@      @      @      @      @                      @      @                      @      T@      4@      T@      0@      (@      $@      �?      @              @      �?       @               @      �?              &@      @      �?      �?      �?                      �?      $@       @      @              @       @      �?       @      �?                       @       @              Q@      @      4@      @      .@      @      ,@              �?      @      �?       @               @      �?                      @      @              H@      �?     �F@              @      �?      @                      �?              @r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ�ޡhG        hNhG        h<Kh=Kh>h"h#K �r�  h%�r�  Rr�  (KK�r�  hV�C              �?r�  tr�  bhJhZhEC       r�  �r�  Rr�  h^Kh_h`Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hE�C       r�  tr�  bK�r�  Rr�  }r�  (hKhjKYhkh"h#K �r�  h%�r�  Rr�  (KKY�r�  hr�Bx         $                   �`@�=����?�             j@                         @�A�d�����?0            @R@������������������������       �                     &@                        p=
�?�^�����?)             O@                         p�A      �?             D@                          @@@     ��?             @@                          �`@X�<ݚ�?             "@������������������������       �                      @	       
       	             �?����X�?             @������������������������       �                      @                          �`@���Q��?             @������������������������       �                     @������������������������       �                      @                           �?�nkK�?             7@������������������������       �        	             .@                        ����?      �?              @                          �`@�q�q�?             @������������������������       �                     �?                         `HA      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                         ��A      �?              @������������������������       �                     @                           @P@      �?             @������������������������       �                     @������������������������       �                     �?       #                   p`@��2(&�?             6@       "                    �P@      �?             @                          �^@      �?             @������������������������       �                      @        !                 ���@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �        
             0@%       X                  ��@������?U             a@&       M                   A�������?T            �`@'       B                   �q@��G���?E            �[@(       A                   �p@��0u���?&             N@)       ,                   �Z@P̏����?%            �L@*       +                   �6@�IєX�?             1@������������������������       �                     �?������������������������       �                     0@-       2                   �
A�G�z�?             D@.       1                  �?A؇���X�?	             ,@/       0                    `P@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     &@3       :                   �;@
j*D>�?             :@4       7       	             �?z�G�z�?             $@5       6                  �&A      �?              @������������������������       �                     �?������������������������       �                     �?8       9                    @K@      �?              @������������������������       �                     �?������������������������       �                     @;       <                     P@     ��?
             0@������������������������       �                     "@=       @                     S@և���X�?             @>       ?                    �?�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?������������������������       �                     @C       L                   ��@�:�]��?            �I@D       K                   H�@PN��T'�?             ;@E       J                  ��AHP�s��?             9@F       I                    �?�q�q�?             @G       H                  �CAz�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �        
             3@������������������������       �                      @������������������������       �                     8@N       Q                  p�A���|���?             6@O       P                 ����?�q�q�?             "@������������������������       �                     @������������������������       �                     @R       S                    9@8�Z$���?	             *@������������������������       �                     �?T       U                    �?�8��8��?             (@������������������������       �                     "@V       W       
             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KKYKK�r�  hV�B�        a@      R@     �@@      D@              &@     �@@      =@      >@      $@      ;@      @      @      @               @      @       @       @              @       @      @                       @      6@      �?      .@              @      �?       @      �?      �?              �?      �?      �?                      �?      @              @      @              @      @      �?      @                      �?      @      3@      @      @      �?      @               @      �?      �?              �?      �?               @                      0@      Z@      @@      Z@      =@     �V@      5@     �E@      1@     �E@      ,@      0@      �?              �?      0@              ;@      *@      (@       @      �?       @      �?                       @      &@              .@      &@       @       @      �?      �?              �?      �?              �?      @      �?                      @      *@      @      "@              @      @      @       @      @                       @              �?              @     �G@      @      7@      @      7@       @      @       @      @      �?      @                      �?              �?      3@                       @      8@              ,@       @      @      @      @                      @      &@       @              �?      &@      �?      "@               @      �?       @                      �?              @r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJQY%hG        hNhG        h<Kh=Kh>h"h#K �r�  h%�r�  Rr�  (KK�r�  hV�C              �?r�  tr�  bhJhZhEC       r�  �r�  Rr�  h^Kh_h`Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hE�C       r�  tr�  bK�r�  Rr�  }r�  (hKhjKUhkh"h#K �r�  h%�r�  Rr�  (KKU�r�  hr�B�                            �`@�����m�?�             j@                           �S@|��?���?#             K@                          �A��V�I��?            �G@������������������������       �                     @                            K@�&!��?            �E@                           �?"pc�
�?             &@                        033�?ףp=
�?             $@������������������������       �                      @	       
                     G@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?                        p=
�?     ��?             @@                           @Q@�KM�]�?             3@������������������������       �                     "@              	             �?z�G�z�?             $@                           �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     *@������������������������       �                     @       L                   �a@tݹ��B�?`            `c@       E                    �Q@lQ���?T            `a@       ,                  �tA�J�4�?L            @_@                        pff�? ,��-�?#            �M@                           �P@�?�|�?            �B@������������������������       �                     @@                           �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?        '                   @@@��2(&�?             6@!       "                   �`@      �?             @������������������������       �                     �?#       $                   �b@�q�q�?             @������������������������       �                     �?%       &                  ��A      �?              @������������������������       �                     �?������������������������       �                     �?(       +                    �?�X�<ݺ?             2@)       *                   �Ar�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     (@-       .                   �;@r٣����?)            �P@������������������������       �                     @/       D                  ��@r�q��?%             N@0       9                    �M@@�r-��?$            �M@1       8                   �C@��p\�?            �D@2       3                 ����?H%u��?             9@������������������������       �                     &@4       5                 �uAd}h���?	             ,@������������������������       �                     @6       7                 pff�?      �?              @������������������������       �                     @������������������������       �                     @������������������������       �        
             0@:       ;                 pff�?�q�q�?             2@������������������������       �                      @<       =                 `ff�?      �?             0@������������������������       �                     "@>       A       	             �?և���X�?             @?       @                 pff�?      �?             @������������������������       �                     @������������������������       �                     �?B       C                   a@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?F       K                  ��A      �?             ,@G       J                 `ff�?�z�G��?             $@H       I                   �f@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @M       R                    �?      �?             0@N       O                 pff�?      �?              @������������������������       �                     @P       Q                   �H@      �?             @������������������������       �                     @������������������������       �                     �?S       T                   @@@      �?              @������������������������       �                     �?������������������������       �                     @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KKUKK�r�  hV�BP        b@     @P@      :@      <@      :@      5@              @      :@      1@      "@       @      "@      �?       @              �?      �?      �?                      �?              �?      1@      .@      1@       @      "@               @       @      �?       @      �?                       @      @                      *@              @     �]@     �B@      \@      ;@     @Z@      4@     �K@      @      B@      �?      @@              @      �?      @                      �?      3@      @       @       @              �?       @      �?      �?              �?      �?      �?                      �?      1@      �?      @      �?      @                      �?      (@              I@      0@              @      I@      $@      I@      "@      C@      @      6@      @      &@              &@      @      @              @      @              @      @              0@              (@      @               @      (@      @      "@              @      @      �?      @              @      �?               @      �?              �?       @                      �?      @      @      @      @      @      �?              �?      @                      @      @              @      $@      @      @      @              �?      @              @      �?              �?      @      �?                      @r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ��fbhG        hNhG        h<Kh=Kh>h"h#K �r�  h%�r�  Rr�  (KK�r�  hV�C              �?r�  tr�  bhJhZhEC       r�  �r�  Rr�  h^Kh_h`Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hE�C       r�  tr�  bK�r�  Rr�  }r�  (hKhjKIhkh"h#K �r�  h%�r�  Rr�  (KKI�r�  hr�B�         (                 p=
�?��Jy(F�?�             j@       	                   �;@j��>��?T            ``@                         P�Ab�2�tk�?
             2@                        ����?"pc�
�?             &@������������������������       �                     "@������������������������       �                      @              
             �?����X�?             @������������������������       �                     @������������������������       �                      @
       '                    `S@hdpZ�L�?J            @\@       $                   �@ ѯ��?G            �Z@                           `@`'�J�?C            �Y@������������������������       �                     �?       #       
             �?T��,��?B            @Y@                          �G@`2U0*��?0            �R@                           �?�O4R���?"            �J@                           �?Pa�	�?            �@@                        `ff�?@4և���?
             ,@������������������������       �                      @                           �?r�q��?             @������������������������       �                     @                         0A      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     3@������������������������       �                     4@       "                   �a@�C��2(�?             6@                        ��A���N8�?             5@������������������������       �                     *@                           �?      �?              @������������������������       �                     @        !                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     :@%       &                  �IA���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @)       *                   �6@$��m��?/            �S@������������������������       �        
             3@+       F                   0�@����*��?%            �M@,       ?                 ���@f�Sc��?            �H@-       6                  @eA�4F����?            �D@.       1                   �A�KM�]�?             3@/       0                   `V@      �?              @������������������������       �                     �?������������������������       �                     �?2       3                   8p@�IєX�?	             1@������������������������       �                     &@4       5                   �G@r�q��?             @������������������������       �                     @������������������������       �                     �?7       >                   `a@      �?             6@8       9                   ��K@D�n�3�?             3@������������������������       �                     @:       ;                    W@������?	             .@������������������������       �                     �?<       =                   �;@d}h���?             ,@������������������������       �                     @������������������������       �                     &@������������������������       �                     @@       A                    O@      �?              @������������������������       �                      @B       C                 ���@r�q��?             @������������������������       �                     @D       E                 033@�q�q�?             @������������������������       �                     �?������������������������       �                      @G       H                   �a@ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KKIKK�r�  hV�B�       �`@     �R@      [@      7@      @      &@       @      "@              "@       @              @       @      @                       @     @Y@      (@     @Y@      @     �X@      @              �?     �X@      @      R@      @      J@      �?      @@      �?      *@      �?       @              @      �?      @              �?      �?      �?                      �?      3@              4@              4@       @      4@      �?      *@              @      �?      @               @      �?       @                      �?              �?      :@              @       @               @      @                      @      ;@     �I@              3@      ;@      @@      2@      ?@      *@      <@       @      1@      �?      �?      �?                      �?      �?      0@              &@      �?      @              @      �?              &@      &@       @      &@      @              @      &@      �?              @      &@      @                      &@      @              @      @               @      @      �?      @               @      �?              �?       @              "@      �?      "@                      �?r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ$�phG        hNhG        h<Kh=Kh>h"h#K �r�  h%�r�  Rr�  (KK�r�  hV�C              �?r�  tr�  bhJhZhEC       r�  �r�  Rr�  h^Kh_h`Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hE�C       r   tr  bK�r  Rr  }r  (hK
hjKYhkh"h#K �r  h%�r  Rr  (KKY�r  hr�Bx                             �`@�����m�?�             j@                           �?�)�8��?)             Q@                         `T	A�Q����?             D@������������������������       �                      @                           @K@     ��?             @@������������������������       �                     "@                          0�@\X��t�?             7@������������������������       �                     "@	                          ґ@����X�?             ,@
                        033�?r�q��?             (@                           �Q@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                      @                           �S@X�Cc�?             <@                          @E@�	j*D�?             :@                          �`@���Q��?             4@                           �H@�z�G��?             $@                          @@@      �?             @              	             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @                          �;@ףp=
�?             $@              
             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @!       6                   @@@��+-l�?b            �a@"       1                  ��A      �?             D@#       0                    �P@��X��?             <@$       '                   �`@�q�q�?             8@%       &                 ���@      �?             @������������������������       �                     @������������������������       �                     �?(       )                    �?ףp=
�?             4@������������������������       �                     $@*       -                    �?z�G�z�?             $@+       ,                   a@      �?              @������������������������       �                     �?������������������������       �                     @.       /                   @k@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @2       3                   d�@�8��8��?             (@������������������������       �                     "@4       5                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @7       V                   �a@�DÓ ��?H            @Y@8       U                  ��@������?D            @X@9       P                   pa@�KM�]�?C            �W@:       G                  P�APN��T'�?'             K@;       B                   @E@��p\�?            �D@<       =                    �? ��WV�?             :@������������������������       �        
             .@>       ?                    �?�C��2(�?
             &@������������������������       �                      @@       A                 ����?�q�q�?             @������������������������       �                      @������������������������       �                     �?C       F                   �G@�r����?
             .@D       E                    �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     $@H       K                    �?�n_Y�K�?	             *@I       J                  0�A      �?              @������������������������       �                      @������������������������       �                     @L       M       
             �?���Q��?             @������������������������       �                     �?N       O                   �D@      �?             @������������������������       �                     @������������������������       �                     �?Q       T                 033@������?            �D@R       S                     T@�(\����?             D@������������������������       �                    �C@������������������������       �                     �?������������������������       �                     �?������������������������       �                      @W       X                    �?      �?             @������������������������       �                      @������������������������       �                      @r	  tr
  bh�h"h#K �r  h%�r  Rr  (KKYKK�r  hV�B�        b@     @P@     �B@      ?@      3@      5@               @      3@      *@      "@              $@      *@              "@      $@      @      $@       @       @       @       @                       @       @                       @      2@      $@      2@       @      (@       @      @      @      @      �?      �?      �?              �?      �?               @                      @      "@      �?       @      �?       @                      �?      @              @                       @     �Z@      A@      4@      4@      3@      "@      3@      @      �?      @              @      �?              2@       @      $@               @       @      @      �?              �?      @              �?      �?      �?                      �?              @      �?      &@              "@      �?       @      �?                       @     �U@      ,@     @U@      (@     @U@      $@      G@       @      C@      @      9@      �?      .@              $@      �?       @               @      �?       @                      �?      *@       @      @       @      @                       @      $@               @      @      @       @               @      @               @      @      �?              �?      @              @      �?             �C@       @     �C@      �?     �C@                      �?              �?               @       @       @       @                       @r  tr  bubhhubh)�r  }r  (hhh	h
hNhKhKhG        hh hNhJW:+LhG        hNhG        h<Kh=Kh>h"h#K �r  h%�r  Rr  (KK�r  hV�C              �?r  tr  bhJhZhEC       r  �r  Rr  h^Kh_h`Kh"h#K �r  h%�r  Rr  (KK�r  hE�C       r   tr!  bK�r"  Rr#  }r$  (hK
hjKQhkh"h#K �r%  h%�r&  Rr'  (KKQ�r(  hr�B�         8                 ����?�����m�?�             j@       1                    �S@f�8A_�?_            �b@                        ����?`����?X            �a@              
             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?       "                  p"A�S</�z�?V            `a@                          �;@h�WH��?A             [@	       
                 `ff�?�n_Y�K�?	             *@������������������������       �                      @                         ��A���!pc�?             &@������������������������       �                      @                           �P@�����H�?             "@������������������������       �                     @              	             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?       !                   ϳ@�}�+r��?8            �W@                          5	A`�q�0ܴ?7            �W@                           �?l��\��?             A@              	             �? ��WV�?             :@                           �?؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     3@                        pff�?      �?              @������������������������       �                     @������������������������       �                      @                         ��A �.�?Ƞ?"             N@������������������������       �                     J@                          P�A      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?#       (                   a@��a�n`�?             ?@$       '                    @P@և���X�?             @%       &                   �B@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @)       ,                   @@@      �?             8@*       +                  �A�q�q�?             @������������������������       �                      @������������������������       �                     @-       0                   �a@�X�<ݺ?             2@.       /                   �[@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �        	             .@2       7                   �`@X�<ݚ�?             "@3       4                    F@r�q��?             @������������������������       �                      @5       6                   <�@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @9       N                    �?����S��?'             M@:       =                    �L@j���� �?             A@;       <                   ��@r�q��?             @������������������������       �                     �?������������������������       �                     @>       ?                   ``@��X��?             <@������������������������       �                     @@       E                  PcA�+e�X�?             9@A       B                    `Q@��S�ۿ?
             .@������������������������       �                     &@C       D                     R@      �?             @������������������������       �                     �?������������������������       �                     @F       G                   �Y@      �?             $@������������������������       �                      @H       K       	             �?      �?              @I       J                 `ff�?�q�q�?             @������������������������       �                     �?������������������������       �                      @L       M                   �*N@���Q��?             @������������������������       �                      @������������������������       �                     @O       P                   �F@      �?             8@������������������������       �                     5@������������������������       �                     @r)  tr*  bh�h"h#K �r+  h%�r,  Rr-  (KKQKK�r.  hV�B        b@     @P@     �_@      8@     �^@      3@      �?       @               @      �?             �^@      1@     �X@      $@       @      @               @       @      @               @       @      �?      @               @      �?       @                      �?     �V@      @     �V@      @      ?@      @      9@      �?      @      �?      @                      �?      3@              @       @      @                       @     �M@      �?      J@              @      �?              �?      @                      �?      8@      @      @      @      @       @               @      @                       @      5@      @      @       @               @      @              1@      �?       @      �?       @                      �?      .@              @      @      �?      @               @      �?      @              @      �?              @              1@     �D@      ,@      4@      @      �?              �?      @              "@      3@      @              @      3@      �?      ,@              &@      �?      @      �?                      @      @      @       @              @      @      �?       @      �?                       @       @      @       @                      @      @      5@              5@      @        r/  tr0  bubhhubh)�r1  }r2  (hhh	h
hNhKhKhG        hh hNhJF<KdhG        hNhG        h<Kh=Kh>h"h#K �r3  h%�r4  Rr5  (KK�r6  hV�C              �?r7  tr8  bhJhZhEC       r9  �r:  Rr;  h^Kh_h`Kh"h#K �r<  h%�r=  Rr>  (KK�r?  hE�C       r@  trA  bK�rB  RrC  }rD  (hK
hjKKhkh"h#K �rE  h%�rF  RrG  (KKK�rH  hr�Bh         *                    �P@6�	���?�             j@                        ����?0z���?_             c@                          �6@�? Da�?N            �_@������������������������       �                     @                          ʶ@�8��8��?I             ^@       	                   0`@؞�z�̼?G            @]@                         ��A      �?             @������������������������       �                     @������������������������       �                     @
                         @�@�v�ɱ?D            �[@                          pa@      �?              @������������������������       �                     �?������������������������       �                     �?              	             �?бK/eh�?B            @[@                         `T	A�}�+r��?             C@                         �9A�q�q�?             @������������������������       �                     �?                           �O@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                    �A@                           �? ��PUp�?'            �Q@������������������������       �                    �I@                           �?P���Q�?             4@������������������������       �        
             1@                           �N@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @       %                   Pr@X�<ݚ�?             ;@                           �M@�<ݚ�?             2@������������������������       �                     @!       $                    �?��S�ۿ?	             .@"       #                     O@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @&       )                    �?�����H�?             "@'       (                 �p=�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @+       @                    �?      �?%             L@,       7                   �`@�ʻ����?             A@-       .                   `@      �?	             0@������������������������       �                      @/       0                  �A����X�?             ,@������������������������       �                     �?1       6                   P�@�θ�?             *@2       5                    @S@�C��2(�?             &@3       4                    �Q@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                      @8       =                   �a@�E��ӭ�?             2@9       :                 ����?8�Z$���?	             *@������������������������       �                     @;       <                    �?�q�q�?             @������������������������       �                      @������������������������       �                     @>       ?                 p=
�?���Q��?             @������������������������       �                      @������������������������       �                     @A       B                   �D@8�A�0��?             6@������������������������       �                     $@C       H                 ��A      �?             (@D       E                    �?�����H�?             "@������������������������       �                     @F       G                   �u@      �?              @������������������������       �                     �?������������������������       �                     �?I       J                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @rI  trJ  bh�h"h#K �rK  h%�rL  RrM  (KKKKK�rN  hV�B�       �b@     �M@     �^@      ?@     �[@      0@              @     �[@      $@     �[@      @      @      @              @      @             �Z@      @      �?      �?      �?                      �?     �Z@      @      B@       @      �?       @              �?      �?      �?              �?      �?             �A@             �Q@      �?     �I@              3@      �?      1@               @      �?              �?       @                      @      (@      .@      @      ,@      @              �?      ,@      �?      @              @      �?                       @       @      �?      �?      �?      �?                      �?      @              <@      <@      3@      .@      @      $@       @              @      $@      �?              @      $@      �?      $@      �?       @               @      �?                       @       @              *@      @      &@       @      @              @       @               @      @               @      @       @                      @      "@      *@              $@      "@      @       @      �?      @              �?      �?      �?                      �?      �?       @      �?                       @rO  trP  bubhhubh)�rQ  }rR  (hhh	h
hNhKhKhG        hh hNhJؽ�hG        hNhG        h<Kh=Kh>h"h#K �rS  h%�rT  RrU  (KK�rV  hV�C              �?rW  trX  bhJhZhEC       rY  �rZ  Rr[  h^Kh_h`Kh"h#K �r\  h%�r]  Rr^  (KK�r_  hE�C       r`  tra  bK�rb  Rrc  }rd  (hKhjK[hkh"h#K �re  h%�rf  Rrg  (KK[�rh  hr�B�                            �`@p�ݯ��?�             j@                          �_@����"�?(             M@������������������������       �                     @                           @K@�b��[��?&            �K@                           1@�q�q�?             .@������������������������       �                      @       
                    y@�θ�?
             *@       	                   jA�q�q�?             @������������������������       �                     �?������������������������       �                      @                         ��Aףp=
�?             $@������������������������       �                     �?������������������������       �                     "@                        ����?R���Q�?             D@������������������������       �                     @                        p=
�?(N:!���?            �A@                        ����?����X�?             ,@                          �`@�θ�?
             *@������������������������       �                     @                          ��@      �?              @                          �a@r�q��?             @������������������������       �                     @              	             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     �?������������������������       �                     5@       T                  �/A�m�tQ�?^            �b@       S                  ��@�'�`d�?Q            �`@       0                    �?z�G�z�?P            @`@        '                   a@�U�=���?*            �P@!       &                  p"Ar�q��?
             2@"       %                   @@@      �?	             0@#       $                    �I@�����H�?             "@������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @(       )                    �P@ �q�q�?              H@������������������������       �                     E@*       /                   �C@�q�q�?             @+       .                   �?@�q�q�?             @,       -                    �R@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @1       @                  @wA     8�?&             P@2       7                   �AX�<ݚ�?             ;@3       4                   `w@ףp=
�?             $@������������������������       �                      @5       6       	             �?      �?              @������������������������       �                     �?������������������������       �                     �?8       =                  @ 
A@�0�!��?             1@9       <                   �a@�r����?             .@:       ;                   h@"pc�
�?             &@������������������������       �                     "@������������������������       �                      @������������������������       �                     @>       ?                    �?      �?              @������������������������       �                     �?������������������������       �                     �?A       R                 �p=�?�MI8d�?            �B@B       C                 033�?�+e�X�?             9@������������������������       �                     @D       M                  0A�q�q�?             2@E       L                   �a@X�<ݚ�?             "@F       G                   �A����X�?             @������������������������       �                     �?H       I                    �?r�q��?             @������������������������       �                     @J       K                 ����?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @N       O                    �?�����H�?             "@������������������������       �                     @P       Q                   @@@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     (@������������������������       �                      @U       X                     J@�����?             3@V       W                   �@����X�?             @������������������������       �                     @������������������������       �                      @Y       Z                   �H@�8��8��?             (@������������������������       �                     &@������������������������       �                     �?ri  trj  bh�h"h#K �rk  h%�rl  Rrm  (KK[KK�rn  hV�B�       �`@     @S@      6@      B@      @              3@      B@      $@      @               @      $@      @      �?       @      �?                       @      "@      �?              �?      "@              "@      ?@      @              @      ?@      @      $@      @      $@              @      @      @      �?      @              @      �?       @      �?                       @       @              �?                      5@     �[@     �D@      Z@      <@      Z@      :@     �N@      @      .@      @      .@      �?       @      �?              �?       @              @                       @      G@       @      E@              @       @      �?       @      �?      �?              �?      �?                      �?      @             �E@      5@      (@      .@      "@      �?       @              �?      �?      �?                      �?      @      ,@       @      *@       @      "@              "@       @                      @      �?      �?      �?                      �?      ?@      @      3@      @      @              (@      @      @      @       @      @      �?              �?      @              @      �?       @      �?                       @       @               @      �?      @              �?      �?              �?      �?              (@                       @      @      *@      @       @      @                       @      �?      &@              &@      �?        ro  trp  bubhhubh)�rq  }rr  (hhh	h
hNhKhKhG        hh hNhJX��vhG        hNhG        h<Kh=Kh>h"h#K �rs  h%�rt  Rru  (KK�rv  hV�C              �?rw  trx  bhJhZhEC       ry  �rz  Rr{  h^Kh_h`Kh"h#K �r|  h%�r}  Rr~  (KK�r  hE�C       r�  tr�  bK�r�  Rr�  }r�  (hKhjKQhkh"h#K �r�  h%�r�  Rr�  (KKQ�r�  hr�B�                 	             �?���֥�?�             j@       	                   �`@���Q��?-            �Q@                           `@��S�ۿ?             .@������������������������       �                     @                           �H@      �?              @                          @@@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @
                            L@^(��I�?%            �K@                         �D�@P���Q�?             4@������������������������       �                     �?������������������������       �                     3@                        `ff�?<=�,S��?            �A@������������������������       �                     @                           �N@���>4��?             <@                         ��A�	j*D�?             *@������������������������       �                      @                          @A"pc�
�?             &@������������������������       �                     @                           �?�q�q�?             @������������������������       �                      @                           �?      �?             @������������������������       �                      @������������������������       �                      @                        fA������?             .@                          �a@      �?              @                           �?�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     @!       "                   �6@�*��?]            `a@������������������������       �                     "@#       >                     Q@
��[��?U            @`@$       /                   �;@�Ra����?<             V@%       .                   N�@�q�q�?             2@&       -                   �q@�t����?             1@'       ,                     P@�q�q�?             (@(       +                   pi@�<ݚ�?             "@)       *                   �b@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     �?0       =       
             �? >�֕�?/            �Q@1       <                 833@��-�=��?            �C@2       ;                    �?�˹�m��?             C@3       :                   ų@z�G�z�?             .@4       5                  ��A؇���X�?
             ,@������������������������       �                     "@6       7                    �?���Q��?             @������������������������       �                      @8       9                   �`@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     7@������������������������       �                     �?������������������������       �                     ?@?       L                   Pa@�ՙ/�?             E@@       A                  `HAl��[B��?             =@������������������������       �                      @B       K                   �`@����X�?             5@C       H                   �G@�t����?             1@D       G                   p`@$�q-�?	             *@E       F                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     $@I       J                   <�@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @M       P                   �?@8�Z$���?             *@N       O                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     "@r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KKQKK�r�  hV�B        a@     @R@      E@      <@      �?      ,@              @      �?      @      �?      @              @      �?                      @     �D@      ,@      3@      �?              �?      3@              6@      *@      @              .@      *@      @      "@       @               @      "@              @       @      @               @       @       @               @       @              &@      @      @      @      @       @               @      @                       @      @             �W@     �F@              "@     �W@      B@     �S@      $@      (@      @      (@      @      @      @      @       @      @       @      @                       @      @                      @      @                      �?     �P@      @     �A@      @     �A@      @      (@      @      (@       @      "@              @       @       @              �?       @      �?                       @              �?      7@                      �?      ?@              0@      :@      ,@      .@       @              @      .@       @      .@      �?      (@      �?       @               @      �?                      $@      �?      @              @      �?              @               @      &@       @       @       @                       @              "@r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ���EhG        hNhG        h<Kh=Kh>h"h#K �r�  h%�r�  Rr�  (KK�r�  hV�C              �?r�  tr�  bhJhZhEC       r�  �r�  Rr�  h^Kh_h`Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hE�C       r�  tr�  bK�r�  Rr�  }r�  (hKhjKOhkh"h#K �r�  h%�r�  Rr�  (KKO�r�  hr�BH                            �6@��+s�?}             j@������������������������       �                     7@       L                    �S@�/�L���?r            @g@       #                   @@@:���١�?k             f@       
                   `@z�):���?             I@                           a@$�q-�?             *@������������������������       �                     "@       	                   �;@      �?             @������������������������       �                     @������������������������       �                     �?                         �OAV������?            �B@                           �P@d}h���?             <@                          �A�LQ�1	�?             7@                         `�
A      �?              @              
             �?r�q��?             @                          0a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �        	             .@                           �Q@���Q��?             @������������������������       �                      @                           �R@�q�q�?             @������������������������       �                      @������������������������       �                     �?                        `ff�?X�<ݚ�?             "@������������������������       �                      @       "                    �M@����X�?             @       !                    @M@r�q��?             @                           ��@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?$       ?                    �?��d��?L            �_@%       :                   �a@Ĝ�oV4�?3            �V@&       /                   �G@ĴF���?-            �T@'       (                   A�i�y�?#            �O@������������������������       �                     >@)       .                   ϳ@�FVQ&�?            �@@*       -                   @A      �?             @@+       ,                   �`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     >@������������������������       �                     �?0       1                   �^@�d�����?
             3@������������������������       �                      @2       9                    �?@�0�!��?	             1@3       4                 ����?�q�q�?             "@������������������������       �                      @5       6                    �?؇���X�?             @������������������������       �                     @7       8                   �K@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @;       <                    �N@X�<ݚ�?             "@������������������������       �                     @=       >                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?@       K                  �A��R[s�?            �A@A       D                 ����?�'�`d�?            �@@B       C                    `@���7�?             6@������������������������       �                     �?������������������������       �                     5@E       J                   �@�eP*L��?             &@F       G                   @B@      �?              @������������������������       �                     �?H       I                    S@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @M       N                  @Aףp=
�?             $@������������������������       �                     �?������������������������       �                     "@r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KKOKK�r�  hV�B�       �`@     �R@              7@     �`@      J@     �`@     �E@      ;@      7@      �?      (@              "@      �?      @              @      �?              :@      &@      6@      @      4@      @      @      @      @      �?      �?      �?              �?      �?              @                       @      .@               @      @               @       @      �?       @                      �?      @      @       @               @      @      �?      @      �?       @      �?                       @              @      �?             �Z@      4@      T@      &@     �R@      @     �N@       @      >@              ?@       @      ?@      �?      �?      �?              �?      �?              >@                      �?      ,@      @               @      ,@      @      @      @               @      @      �?      @               @      �?       @                      �?       @              @      @              @      @      �?      @                      �?      :@      "@      :@      @      5@      �?              �?      5@              @      @       @      @      �?              �?      @      �?                      @      @                       @      �?      "@      �?                      "@r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ:9)bhG        hNhG        h<Kh=Kh>h"h#K �r�  h%�r�  Rr�  (KK�r�  hV�C              �?r�  tr�  bhJhZhEC       r�  �r�  Rr�  h^Kh_h`Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hE�C       r�  tr�  bK�r�  Rr�  }r�  (hKhjKMhkh"h#K �r�  h%�r�  Rr�  (KKM�r�  hr�B�                            �6@�oUN�1�?}             j@������������������������       �                     8@       (                   �`@���@��?r             g@                           �?��k��?$            �J@                          �C@���|���?            �@@                           w@      �?             4@       
                  `T	A���!pc�?             &@       	                 pff�?      �?              @������������������������       �                     �?������������������������       �                     @                            P@�q�q�?             @������������������������       �                      @������������������������       �                     �?              	             �?�<ݚ�?             "@                          �`@      �?              @������������������������       �                     �?������������������������       �                     �?                         ��A؇���X�?             @������������������������       �                     �?������������������������       �                     @                          �^@8�Z$���?	             *@������������������������       �                     �?              	             �?�8��8��?             (@������������������������       �                     @                          �K@؇���X�?             @������������������������       �                     @������������������������       �                     �?       #                    �?���Q��?             4@                           �?      �?              @������������������������       �                     @       "       
             �?���Q��?             @        !                   �`@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?$       %                   d	A      �?             (@������������������������       �                      @&       '                   X@ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?)       .                 033�?<���D�?N            �`@*       +                    �?XB���?             =@������������������������       �                     2@,       -                  �A�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?/       H                     S@�	��)��?;            �Y@0       3                  @�@�¦�{��?7            �W@1       2                   Ȗ@      �?              @������������������������       �                     �?������������������������       �                     �?4       ;                  ��A��y� �?5            @W@5       :                    @J@@��8��?             H@6       9                   a@      �?             0@7       8       
             �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     &@������������������������       �                     @@<       G                 �p=�?���V��?            �F@=       >                 `ff�?8����?             7@������������������������       �                     @?       F                   �C@j���� �?             1@@       E                   �@��
ц��?	             *@A       B                    �?�q�q�?             "@������������������������       �                     @C       D                   �W@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �        	             6@I       L                    �?      �?              @J       K       
             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KKMKK�r�  hV�B�        b@      P@              8@      b@      D@      =@      8@      5@      (@      $@      $@      @       @      �?      @      �?                      @       @      �?       @                      �?      @       @      �?      �?      �?                      �?      @      �?              �?      @              &@       @              �?      &@      �?      @              @      �?      @                      �?       @      (@      @      @      @               @      @      �?      @      �?                      @      �?              @      "@       @              �?      "@              "@      �?              ]@      0@      <@      �?      2@              $@      �?      $@                      �?      V@      .@     �U@      "@      �?      �?      �?                      �?     @U@       @     �G@      �?      .@      �?      @      �?      @                      �?      &@              @@              C@      @      0@      @      @              $@      @      @      @      @      @      @              �?      @      �?                      @              @      @              6@               @      @       @      �?       @                      �?              @r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ�BHzhG        hNhG        h<Kh=Kh>h"h#K �r�  h%�r�  Rr�  (KK�r�  hV�C              �?r�  tr�  bhJhZhEC       r�  �r�  Rr�  h^Kh_h`Kh"h#K �r�  h%�r�  Rr�  (KK�r�  hE�C       r�  tr�  bK�r�  Rr�  }r�  (hKhjKIhkh"h#K �r�  h%�r�  Rr�  (KKI�r�  hr�B�                             @@@��+s�?�             j@                          �`@     ��?&             P@                        ����?`2U0*��?             9@                          ��@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     6@                           �?��Zy�?            �C@	                          ��@      �?             0@
                        ����?����X�?             ,@������������������������       �                     @                          �V@և���X�?             @������������������������       �                     �?              
             �?�q�q�?             @������������������������       �                      @                           �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @                          �a@8����?             7@                           @O@�S����?             3@              
             �?      �?             (@                          @A      �?             @������������������������       �                     �?                           �?�q�q�?             @������������������������       �                     �?������������������������       �                      @                         @�A      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @!       B                    �S@z�G�z�?b             b@"       =                 ����?X�EQ]N�?X             `@#       0                     Q@T(y2��?P            �]@$       +                   �a@x��B�R�?@            �V@%       &                  p"A �)���?8            @T@������������������������       �        ,             P@'       (                    �?�IєX�?             1@������������������������       �        
             .@)       *                 ����?      �?              @������������������������       �                     �?������������������������       �                     �?,       -                    �@z�G�z�?             $@������������������������       �                     @.       /                  8�A�q�q�?             @������������������������       �                      @������������������������       �                     �?1       6                    �?�>4և��?             <@2       3                   @J@      �?	             0@������������������������       �                     &@4       5                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @7       8                   @E@�q�q�?             (@������������������������       �                     @9       <       
             �?և���X�?             @:       ;                   �X@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @>       A                 033@�z�G��?             $@?       @                   �S@      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                      @C       D                   �`@      �?
             0@������������������������       �                     (@E       H                    �?      �?             @F       G                 `ff�?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KKIKK�r�  hV�B�       �`@     �R@      2@      G@      �?      8@      �?       @      �?                       @              6@      1@      6@      $@      @      $@      @      @              @      @      �?               @      @               @       @       @       @                       @               @      @      0@      @      0@      @      "@       @       @              �?       @      �?              �?       @              �?      @      �?                      @              @      @              ]@      =@     �\@      .@     �[@       @      V@      @      T@      �?      P@              0@      �?      .@              �?      �?      �?                      �?       @       @      @              �?       @               @      �?              7@      @      .@      �?      &@              @      �?              �?      @               @      @      @              @      @      @       @               @      @                       @      @      @      �?      @      �?                      @       @               @      ,@              (@       @       @      �?       @      �?                       @      �?        r�  tr�  bubhhubehhub.